magic
tech sky130A
magscale 1 2
timestamp 1770916899
<< nwell >>
rect 5398 469 5582 480
rect 3221 41 3341 225
<< pwell >>
rect 2265 -1059 2347 -917
<< viali >>
rect 828 482 959 527
rect 3096 484 3221 530
rect 5426 484 5551 530
rect 2128 -1270 2246 -1220
rect 5425 -1790 5539 -1736
rect 2113 -2629 2236 -2580
<< metal1 >>
rect -584 982 7505 1225
rect 384 221 554 982
rect 804 527 982 982
rect 804 482 828 527
rect 959 482 982 527
rect 804 473 982 482
rect 865 377 1245 424
rect 384 51 876 221
rect 914 51 977 221
rect 1147 51 1153 221
rect 1198 -102 1245 377
rect 2673 229 2857 982
rect 3067 530 3250 982
rect 3067 484 3096 530
rect 3221 484 3250 530
rect 3067 478 3250 484
rect 3128 381 3501 428
rect 2673 45 3138 229
rect 3175 196 3295 229
rect 3169 76 3175 196
rect 3295 76 3301 196
rect 3175 45 3295 76
rect 3454 -98 3501 381
rect 4981 218 5166 982
rect 5398 530 5582 982
rect 5398 484 5426 530
rect 5551 484 5582 530
rect 5398 469 5582 484
rect 6247 436 6304 442
rect 5462 382 6247 427
rect 5462 379 5909 382
rect 6247 372 6304 378
rect 4981 33 5470 218
rect 5508 194 5910 220
rect 5508 69 5759 194
rect 5884 69 5910 194
rect 5508 43 5910 69
rect 3448 -99 3501 -98
rect 6255 -99 6303 372
rect 1197 -103 1245 -102
rect 865 -150 1245 -103
rect 3125 -146 3501 -99
rect 103 -708 303 -663
rect 1197 -708 1244 -150
rect 103 -808 1244 -708
rect 1835 -808 2215 -806
rect 103 -817 2215 -808
rect 103 -863 303 -817
rect 1194 -854 2215 -817
rect 1194 -855 1883 -854
rect 1645 -953 1713 -947
rect 1645 -1354 1713 -1021
rect 1835 -1116 1883 -855
rect 2014 -1052 2020 -922
rect 2150 -1052 2161 -922
rect 2199 -1059 2205 -917
rect 2347 -1059 2353 -917
rect 2207 -1060 2298 -1059
rect 1835 -1164 2213 -1116
rect 2098 -1220 2272 -1210
rect 2098 -1270 2128 -1220
rect 2246 -1270 2272 -1220
rect 2098 -1354 2272 -1270
rect 1645 -1422 2272 -1354
rect 104 -1921 633 -1721
rect 833 -1921 839 -1721
rect 1645 -1843 1713 -1422
rect 2028 -1573 2034 -1521
rect 2086 -1524 2092 -1521
rect 3448 -1524 3495 -146
rect 5461 -147 6303 -99
rect 6250 -1323 6303 -147
rect 6653 -597 6778 -591
rect 7401 -597 7601 -558
rect 6778 -722 7601 -597
rect 6653 -728 6778 -722
rect 7401 -758 7601 -722
rect 5452 -1376 6303 -1323
rect 2086 -1571 3495 -1524
rect 4973 -1568 5464 -1445
rect 2086 -1573 2092 -1571
rect 1645 -1911 2551 -1843
rect 1447 -2166 1499 -2160
rect 1767 -2168 2208 -2167
rect 1499 -2215 2208 -2168
rect 1447 -2224 1499 -2218
rect 1541 -2313 1619 -2307
rect 1541 -2869 1619 -2391
rect 1765 -2478 1813 -2215
rect 2483 -2291 2551 -1911
rect 2026 -2292 2032 -2291
rect 1993 -2413 2032 -2292
rect 2154 -2413 2160 -2291
rect 2198 -2412 2551 -2291
rect 1765 -2526 2206 -2478
rect 2085 -2580 2271 -2566
rect 2085 -2629 2113 -2580
rect 2236 -2629 2271 -2580
rect 2085 -2869 2271 -2629
rect 4973 -2869 5096 -1568
rect 5501 -1569 5759 -1444
rect 5884 -1569 5890 -1444
rect 6250 -1635 6303 -1376
rect 5451 -1688 6303 -1635
rect 5383 -1736 5569 -1729
rect 5383 -1790 5425 -1736
rect 5539 -1790 5569 -1736
rect 5383 -2869 5569 -1790
rect -587 -3132 7509 -2869
<< via1 >>
rect 977 51 1147 221
rect 3175 76 3295 196
rect 6247 378 6304 436
rect 5759 69 5884 194
rect 1645 -1021 1713 -953
rect 2020 -1052 2150 -922
rect 2205 -1059 2347 -917
rect 633 -1921 833 -1721
rect 2034 -1573 2086 -1521
rect 6653 -722 6778 -597
rect 1447 -2218 1499 -2166
rect 1541 -2391 1619 -2313
rect 2032 -2413 2154 -2291
rect 5759 -1569 5884 -1444
<< metal2 >>
rect 1856 724 6305 781
rect 977 221 1147 227
rect 1856 165 1913 724
rect 3633 723 6305 724
rect 3175 196 3295 202
rect 1147 108 1914 165
rect 977 45 1147 51
rect 1860 -491 1914 108
rect 3850 162 3908 723
rect 6247 436 6305 723
rect 6241 378 6247 436
rect 6304 378 6310 436
rect 3295 110 3908 162
rect 5759 194 5884 200
rect 3175 70 3295 76
rect 1860 -558 2647 -491
rect 2020 -922 2150 -916
rect 1639 -1021 1645 -953
rect 1713 -1021 2020 -953
rect 2020 -1058 2150 -1052
rect 2205 -917 2347 -911
rect 2580 -954 2647 -558
rect 2347 -1021 2647 -954
rect 5759 -597 5884 69
rect 5759 -722 6653 -597
rect 6778 -722 6784 -597
rect 2205 -1065 2347 -1059
rect 5759 -1444 5884 -722
rect 2034 -1521 2086 -1515
rect 1449 -1570 2034 -1523
rect 633 -1721 833 -1715
rect 1449 -1788 1496 -1570
rect 2034 -1579 2086 -1573
rect 5759 -1575 5884 -1569
rect 833 -1853 1496 -1788
rect 633 -1927 833 -1921
rect 1449 -2166 1496 -1853
rect 1441 -2218 1447 -2166
rect 1499 -2218 1505 -2166
rect 2032 -2291 2154 -2285
rect 1535 -2391 1541 -2313
rect 1619 -2391 2032 -2313
rect 2032 -2419 2154 -2413
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1770916899
transform 1 0 2181 0 1 -988
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGAKDL  XM2
timestamp 1770916899
transform 1 0 895 0 1 137
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM3
timestamp 1770916899
transform 1 0 3155 0 1 141
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1770916899
transform 1 0 2175 0 1 -2346
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGAKDL  XM5
timestamp 1770916899
transform 1 0 5491 0 1 139
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_648S5X  XM6
timestamp 1770916899
transform 1 0 5481 0 1 -1506
box -211 -310 211 310
<< labels >>
flabel metal1 -495 999 -295 1199 0 FreeSans 256 0 0 0 VCC
port 3 nsew
flabel metal1 -491 -3100 -291 -2900 0 FreeSans 256 0 0 0 GND
port 4 nsew
flabel metal1 104 -1921 304 -1721 0 FreeSans 256 0 0 0 B
port 1 nsew
flabel metal1 103 -863 303 -663 0 FreeSans 256 0 0 0 A
port 0 nsew
flabel metal1 7401 -758 7601 -558 0 FreeSans 256 0 0 0 Y
port 2 nsew
<< end >>
