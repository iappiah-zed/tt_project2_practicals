** sch_path: /home/iappiah/tt_project2_practicals/xschem/AND_IC_TopLevel.sch
.subckt AND_IC_TopLevel 1A 1B 1Y 2A 2B 2Y GND 3A 3B 3Y 4A 4B 4Y VCC
*.PININFO 1A:I GND:B 1Y:O 1B:I 2A:I 2B:I 3A:I 3B:I 4A:I 4B:I 2Y:O 3Y:O 4Y:O VCC:B
x1 1A 1B 1Y VCC GND ic_7804_AND
x2 2A 2B 2Y VCC GND ic_7804_AND
x3 3A 3B 3Y VCC GND ic_7804_AND
x4 4A 4B 4Y VCC GND ic_7804_AND
.ends

* expanding   symbol:  ic_7804_AND.sym # of pins=5
** sym_path: /home/iappiah/tt_project2_practicals/xschem/ic_7804_AND.sym
** sch_path: /home/iappiah/tt_project2_practicals/xschem/ic_7804_AND.sch
.subckt ic_7804_AND A B Y VCC GND
*.PININFO A:I Y:O B:I VCC:B GND:B
XM2 net1 A VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM3 net1 B VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM5 Y net1 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM1 net1 A net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net2 B GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 Y net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
