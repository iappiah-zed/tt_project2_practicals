magic
tech sky130A
magscale 1 2
timestamp 1771576399
<< metal1 >>
rect 1437 33750 1637 33756
rect 1437 33126 1637 33550
rect 19896 31406 19956 31412
rect 6612 31248 6618 31308
rect 6678 31248 6684 31308
rect 7344 31262 7350 31322
rect 7410 31262 7416 31322
rect 4570 31206 4630 31212
rect 4570 21606 4630 31146
rect 5644 30752 5704 30758
rect 5644 22660 5704 30692
rect 6618 29128 6678 31248
rect 7350 30140 7410 31262
rect 16494 31160 16500 31220
rect 16560 31160 16566 31220
rect 16500 30214 16560 31160
rect 19896 30222 19956 31346
rect 28376 30904 28382 30964
rect 28442 30904 28448 30964
rect 28382 30138 28442 30904
rect 28872 29510 28878 29570
rect 28938 29510 28944 29570
rect 6618 29068 7390 29128
rect 28878 29038 28938 29510
rect 29705 25860 30342 26060
rect 28472 23228 28532 23234
rect 28532 23168 29076 23228
rect 28472 23162 28532 23168
rect 19890 22812 19896 22872
rect 19956 22812 19962 22872
rect 5644 22600 7366 22660
rect 16484 22094 16490 22154
rect 16550 22094 16556 22154
rect 4570 21546 7408 21606
rect 16490 21444 16550 22094
rect 19896 21476 19956 22812
rect 29016 22588 29076 23168
rect 29612 21908 29672 21914
rect 29612 21590 29672 21848
rect 29028 21530 29672 21590
rect 30142 21292 30342 25860
rect 30142 21086 30342 21092
<< via1 >>
rect 1437 33550 1637 33750
rect 19896 31346 19956 31406
rect 6618 31248 6678 31308
rect 7350 31262 7410 31322
rect 4570 31146 4630 31206
rect 5644 30692 5704 30752
rect 16500 31160 16560 31220
rect 28382 30904 28442 30964
rect 28878 29510 28938 29570
rect 28472 23168 28532 23228
rect 19896 22812 19956 22872
rect 16490 22094 16550 22154
rect 29612 21848 29672 21908
rect 30142 21092 30342 21292
<< metal2 >>
rect 15166 42720 15222 42727
rect 24344 42720 24404 42729
rect 15164 42718 24344 42720
rect 15164 42662 15166 42718
rect 15222 42662 24344 42718
rect 15164 42660 24344 42662
rect 15166 42653 15222 42660
rect 24344 42651 24404 42660
rect 14040 41812 23798 41872
rect 23858 41812 23867 41872
rect 14040 37676 14100 41812
rect 27116 41602 27176 41611
rect 5644 37616 14100 37676
rect 15164 41184 15224 41193
rect 5058 36754 5118 36763
rect 4570 36694 5058 36754
rect 1437 34164 1637 34173
rect 1437 33750 1637 33964
rect 1431 33550 1437 33750
rect 1637 33550 1643 33750
rect 4570 31206 4630 36694
rect 5058 36685 5118 36694
rect 4564 31146 4570 31206
rect 4630 31146 4636 31206
rect 5644 30752 5704 37616
rect 6208 36754 6264 36761
rect 15164 36754 15224 41124
rect 18832 39196 18892 39205
rect 6206 36752 15224 36754
rect 6206 36696 6208 36752
rect 6264 36696 15224 36752
rect 16500 39136 18832 39196
rect 16500 36726 16560 39136
rect 18832 39127 18892 39136
rect 17172 38524 17232 38533
rect 6206 36694 15224 36696
rect 6208 36687 6264 36694
rect 16493 36670 16502 36726
rect 16558 36670 16567 36726
rect 16500 36668 16560 36670
rect 17172 36586 17232 38464
rect 17165 36530 17174 36586
rect 17230 36530 17239 36586
rect 17172 36528 17232 36530
rect 27116 35846 27176 41542
rect 6618 35786 27176 35846
rect 27660 40574 27720 40583
rect 6618 31308 6678 35786
rect 27660 34972 27720 40514
rect 7350 34912 27720 34972
rect 7350 31322 7410 34912
rect 19887 34330 19896 34390
rect 19956 34330 19965 34390
rect 17172 34302 17232 34311
rect 7350 31256 7410 31262
rect 16500 33968 16560 33977
rect 6618 31242 6678 31248
rect 16500 31220 16560 33908
rect 16500 31154 16560 31160
rect 5638 30692 5644 30752
rect 5704 30692 5710 30752
rect 17172 29158 17232 34242
rect 16490 29098 17232 29158
rect 18212 33934 18272 33943
rect 18212 29158 18272 33874
rect 19896 31406 19956 34330
rect 26004 34290 26064 34299
rect 26064 34230 28938 34290
rect 26004 34221 26064 34230
rect 24282 33632 24342 33641
rect 20972 33572 24282 33632
rect 19890 31346 19896 31406
rect 19956 31346 19962 31406
rect 18212 29098 19956 29158
rect 16490 22154 16550 29098
rect 19896 22872 19956 29098
rect 20972 26242 21032 33572
rect 24282 33563 24342 33572
rect 28382 31254 28442 31256
rect 28375 31198 28384 31254
rect 28440 31198 28449 31254
rect 28382 30964 28442 31198
rect 28382 30898 28442 30904
rect 23996 30832 24056 30841
rect 23996 26904 24056 30772
rect 28878 29570 28938 34230
rect 28878 29504 28938 29510
rect 23996 26844 28134 26904
rect 20972 26182 27440 26242
rect 27380 23228 27440 26182
rect 28074 25232 28134 26844
rect 29612 25232 29672 25236
rect 28074 25172 29672 25232
rect 27380 23168 28472 23228
rect 28532 23168 28538 23228
rect 19896 22806 19956 22812
rect 16490 22088 16550 22094
rect 29612 21908 29672 25172
rect 29606 21848 29612 21908
rect 29672 21848 29678 21908
rect 30136 21092 30142 21292
rect 30342 21092 30348 21292
rect 30142 20230 30342 21092
rect 30142 20021 30342 20030
<< via2 >>
rect 15166 42662 15222 42718
rect 24344 42660 24404 42720
rect 23798 41812 23858 41872
rect 27116 41542 27176 41602
rect 15164 41124 15224 41184
rect 5058 36694 5118 36754
rect 1437 33964 1637 34164
rect 6208 36696 6264 36752
rect 18832 39136 18892 39196
rect 17172 38464 17232 38524
rect 16502 36670 16558 36726
rect 17174 36530 17230 36586
rect 27660 40514 27720 40574
rect 19896 34330 19956 34390
rect 17172 34242 17232 34302
rect 16500 33908 16560 33968
rect 18212 33874 18272 33934
rect 26004 34230 26064 34290
rect 24282 33572 24342 33632
rect 28384 31198 28440 31254
rect 23996 30772 24056 30832
rect 30142 20030 30342 20230
<< metal3 >>
rect 18270 44086 18276 44150
rect 18340 44148 18346 44150
rect 19888 44148 19894 44150
rect 18340 44088 19894 44148
rect 18340 44086 18346 44088
rect 19888 44086 19894 44088
rect 19958 44086 19964 44150
rect 24342 43884 24406 43890
rect 24342 43814 24406 43820
rect 23788 43256 23794 43320
rect 23858 43256 23864 43320
rect 15161 42718 15227 42723
rect 15161 42662 15166 42718
rect 15222 42662 15227 42718
rect 15161 42657 15227 42662
rect 15164 41189 15224 42657
rect 23796 42430 23856 43256
rect 24344 42725 24404 43814
rect 27106 43006 27170 43012
rect 27106 42936 27170 42942
rect 24339 42720 24409 42725
rect 24339 42660 24344 42720
rect 24404 42660 24409 42720
rect 24339 42655 24409 42660
rect 23796 42180 23858 42430
rect 23798 41877 23858 42180
rect 27108 42038 27168 42936
rect 27656 42366 27720 42372
rect 27656 42296 27720 42302
rect 23793 41872 23863 41877
rect 23793 41812 23798 41872
rect 23858 41812 23863 41872
rect 23793 41807 23863 41812
rect 27108 41764 27176 42038
rect 27116 41607 27176 41764
rect 27111 41602 27181 41607
rect 27111 41542 27116 41602
rect 27176 41542 27181 41602
rect 27111 41537 27181 41542
rect 15159 41184 15229 41189
rect 15159 41124 15164 41184
rect 15224 41124 15229 41184
rect 15159 41119 15229 41124
rect 27658 40846 27718 42296
rect 27658 40658 27720 40846
rect 27660 40579 27720 40658
rect 27655 40574 27725 40579
rect 27655 40514 27660 40574
rect 27720 40514 27725 40574
rect 27655 40509 27725 40514
rect 18830 40468 18894 40474
rect 18830 40398 18894 40404
rect 17166 40148 17172 40212
rect 17236 40148 17242 40212
rect 18204 40176 18268 40182
rect 17174 39188 17234 40148
rect 18204 40106 18268 40112
rect 17172 38850 17234 39188
rect 18206 39074 18266 40106
rect 18832 39201 18892 40398
rect 18827 39196 18897 39201
rect 18827 39136 18832 39196
rect 18892 39136 18897 39196
rect 18827 39131 18897 39136
rect 18206 38934 18272 39074
rect 17172 38529 17232 38850
rect 17167 38524 17237 38529
rect 17167 38464 17172 38524
rect 17232 38464 17237 38524
rect 17167 38459 17237 38464
rect 5053 36754 5123 36759
rect 6203 36754 6269 36757
rect 5053 36694 5058 36754
rect 5118 36752 6269 36754
rect 5118 36696 6208 36752
rect 6264 36696 6269 36752
rect 5118 36694 6269 36696
rect 5053 36689 5123 36694
rect 6203 36691 6269 36694
rect 16497 36726 16563 36731
rect 16497 36670 16502 36726
rect 16558 36670 16563 36726
rect 16497 36665 16563 36670
rect 244 34536 250 34736
rect 450 34536 1637 34736
rect 1437 34169 1637 34536
rect 1432 34164 1642 34169
rect 1432 33964 1437 34164
rect 1637 33964 1642 34164
rect 16500 33973 16560 36665
rect 17169 36586 17235 36591
rect 17169 36530 17174 36586
rect 17230 36530 17235 36586
rect 17169 36525 17235 36530
rect 17172 34307 17232 36525
rect 17167 34302 17237 34307
rect 17167 34242 17172 34302
rect 17232 34242 17237 34302
rect 17167 34237 17237 34242
rect 1432 33959 1642 33964
rect 16495 33968 16565 33973
rect 16495 33908 16500 33968
rect 16560 33908 16565 33968
rect 18212 33939 18272 38934
rect 26002 36468 26066 36474
rect 19894 36406 19958 36412
rect 26002 36398 26066 36404
rect 19894 36336 19958 36342
rect 19896 34395 19956 36336
rect 19891 34390 19961 34395
rect 19891 34330 19896 34390
rect 19956 34330 19961 34390
rect 19891 34325 19961 34330
rect 26004 34295 26064 36398
rect 25999 34290 26069 34295
rect 25999 34230 26004 34290
rect 26064 34230 26069 34290
rect 25999 34225 26069 34230
rect 16495 33903 16565 33908
rect 18207 33934 18277 33939
rect 18207 33874 18212 33934
rect 18272 33874 18277 33934
rect 18207 33869 18277 33874
rect 24277 33632 24347 33637
rect 24896 33632 24902 33634
rect 24277 33572 24282 33632
rect 24342 33572 24902 33632
rect 24277 33567 24347 33572
rect 24896 33570 24902 33572
rect 24966 33570 24972 33634
rect 25452 33470 25516 33476
rect 25452 33400 25516 33406
rect 25454 32910 25514 33400
rect 23996 32850 25514 32910
rect 23996 30837 24056 32850
rect 28374 31492 28380 31556
rect 28444 31492 28450 31556
rect 28382 31259 28442 31492
rect 28379 31254 28445 31259
rect 28379 31198 28384 31254
rect 28440 31198 28445 31254
rect 28379 31193 28445 31198
rect 23991 30832 24061 30837
rect 23991 30772 23996 30832
rect 24056 30772 24061 30832
rect 23991 30767 24061 30772
rect 30137 20230 30347 20235
rect 30137 20030 30142 20230
rect 30342 20030 30347 20230
rect 30137 20025 30347 20030
rect 30142 17936 30342 20025
rect 30142 17730 30342 17736
<< via3 >>
rect 18276 44086 18340 44150
rect 19894 44086 19958 44150
rect 24342 43820 24406 43884
rect 23794 43256 23858 43320
rect 27106 42942 27170 43006
rect 27656 42302 27720 42366
rect 18830 40404 18894 40468
rect 17172 40148 17236 40212
rect 18204 40112 18268 40176
rect 250 34536 450 34736
rect 19894 36342 19958 36406
rect 26002 36404 26066 36468
rect 24902 33570 24966 33634
rect 25452 33406 25516 33470
rect 28380 31492 28444 31556
rect 30142 17736 30342 17936
<< metal4 >>
rect 6134 44754 6194 45152
rect 6686 44754 6746 45152
rect 7238 44754 7298 45152
rect 7790 44754 7850 45152
rect 8342 44754 8402 45152
rect 8894 44754 8954 45152
rect 9446 44754 9506 45152
rect 9998 44754 10058 45152
rect 10550 44754 10610 45152
rect 11102 44754 11162 45152
rect 11654 44754 11714 45152
rect 12206 44754 12266 45152
rect 12758 44754 12818 45152
rect 13310 44754 13370 45152
rect 13862 44754 13922 45152
rect 14414 44754 14474 45152
rect 14966 44754 15026 45152
rect 15518 44754 15578 45152
rect 16070 44754 16130 45152
rect 16622 44754 16682 45152
rect 6118 44674 16682 44754
rect 6118 44672 16673 44674
rect 200 34736 600 44152
rect 200 34536 250 34736
rect 450 34536 600 34736
rect 200 1000 600 34536
rect 800 43971 1200 44152
rect 6118 43971 6200 44672
rect 8894 44670 8954 44672
rect 14414 44670 14474 44672
rect 800 43889 6200 43971
rect 800 18026 1200 43889
rect 17174 40213 17234 45152
rect 17726 41092 17786 45152
rect 18278 44151 18338 45152
rect 18275 44150 18341 44151
rect 18275 44086 18276 44150
rect 18340 44086 18341 44150
rect 18275 44085 18341 44086
rect 17726 41032 18266 41092
rect 17171 40212 17237 40213
rect 17171 40148 17172 40212
rect 17236 40148 17237 40212
rect 18206 40177 18266 41032
rect 18830 40770 18890 45152
rect 19382 44950 19442 45152
rect 19934 44950 19994 45152
rect 20486 44950 20546 45152
rect 21038 44950 21098 45152
rect 21590 44950 21650 45152
rect 22142 44950 22202 45152
rect 22694 44950 22754 45152
rect 23246 44950 23306 45152
rect 23798 44582 23858 45152
rect 23796 44454 23858 44582
rect 19893 44150 19959 44151
rect 19893 44086 19894 44150
rect 19958 44086 19959 44150
rect 19893 44085 19959 44086
rect 18830 40596 18892 40770
rect 18832 40469 18892 40596
rect 18829 40468 18895 40469
rect 18829 40404 18830 40468
rect 18894 40404 18895 40468
rect 18829 40403 18895 40404
rect 17171 40147 17237 40148
rect 18203 40176 18269 40177
rect 18203 40112 18204 40176
rect 18268 40112 18269 40176
rect 18203 40111 18269 40112
rect 19896 36407 19956 44085
rect 23796 43321 23856 44454
rect 24350 44364 24410 45152
rect 24348 44222 24410 44364
rect 24348 44162 24408 44222
rect 24344 43980 24408 44162
rect 24344 43885 24404 43980
rect 24341 43884 24407 43885
rect 24341 43820 24342 43884
rect 24406 43820 24407 43884
rect 24341 43819 24407 43820
rect 23793 43320 23859 43321
rect 23793 43256 23794 43320
rect 23858 43256 23859 43320
rect 23793 43255 23859 43256
rect 19893 36406 19959 36407
rect 19893 36342 19894 36406
rect 19958 36342 19959 36406
rect 19893 36341 19959 36342
rect 24902 34344 24962 45152
rect 24902 34244 24964 34344
rect 24904 33635 24964 34244
rect 24901 33634 24967 33635
rect 24901 33570 24902 33634
rect 24966 33570 24967 33634
rect 24901 33569 24967 33570
rect 25454 33471 25514 45152
rect 26006 44463 26066 45152
rect 25985 41003 26071 44463
rect 25998 37148 26058 41003
rect 25998 36812 26064 37148
rect 26004 36469 26064 36812
rect 26001 36468 26067 36469
rect 26001 36404 26002 36468
rect 26066 36404 26067 36468
rect 26001 36403 26067 36404
rect 25451 33470 25517 33471
rect 25451 33406 25452 33470
rect 25516 33406 25517 33470
rect 25451 33405 25517 33406
rect 26558 32894 26618 45152
rect 27110 43488 27170 45152
rect 27108 43254 27170 43488
rect 27108 43007 27168 43254
rect 27105 43006 27171 43007
rect 27105 42942 27106 43006
rect 27170 42942 27171 43006
rect 27662 42984 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27105 42941 27171 42942
rect 27658 42524 27722 42984
rect 27658 42367 27718 42524
rect 27655 42366 27721 42367
rect 27655 42302 27656 42366
rect 27720 42302 27721 42366
rect 27655 42301 27721 42302
rect 26558 32834 28442 32894
rect 28382 31557 28442 32834
rect 28379 31556 28445 31557
rect 28379 31492 28380 31556
rect 28444 31492 28445 31556
rect 28379 31491 28445 31492
rect 800 17936 29072 18026
rect 30141 17936 30343 17937
rect 800 17736 30142 17936
rect 30342 17736 30343 17936
rect 800 17626 29072 17736
rect 30141 17735 30343 17736
rect 800 1000 1200 17626
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use AND_IC_TopLevel  AND_IC_TopLevel_0
timestamp 1771336497
transform 1 0 7561 0 1 33012
box -6143 -13442 22344 346
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
