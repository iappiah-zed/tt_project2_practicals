** sch_path: /home/iappiah/tt_project2_practicals/xschem/AND_IC_TopLevel.sch
.subckt AND_IC_TopLevel 1A 1B 1Y 2A 2B 2Y GND 3A 3B 3Y 4A 4B 4Y VCC
*.PININFO 1A:I GND:B 1Y:O 1B:I 2A:I 2B:I 3A:I 3B:I 4A:I 4B:I 2Y:O 3Y:O 4Y:O VCC:B
x1 1A 1B 1Y VCC GND 7804_AND_IC
x2 2A 2B 2Y VCC GND 7804_AND_IC
x3 3A 3B 3Y VCC GND 7804_AND_IC
x4 4A 4B 4Y VCC GND 7804_AND_IC
D1 1A VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D2 GND 1A sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D3 1B VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D4 GND 1B sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D5 1Y VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D6 GND 1Y sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D7 2Y VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D8 GND 2Y sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D9 2A VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D10 GND 2A sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D11 2B VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D12 GND 2B sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D13 4B VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D14 GND 4B sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D15 4A VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D16 GND 4A sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D17 3A VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D18 GND 3A sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D19 3B VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D20 GND 3B sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D21 4Y VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D22 GND 4Y sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D23 3Y VCC sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D24 GND 3Y sky130_fd_pr__diode_pw2nd_05v5 area=1e12 pj=4e6
D25 GND VCC sky130_fd_pr__diode_pw2nd_05v5 area=100e12 pj=400e6
.ends

* expanding   symbol:  7804_AND_IC.sym # of pins=5
** sym_path: /home/iappiah/tt_project2_practicals/xschem/7804_AND_IC.sym
** sch_path: /home/iappiah/tt_project2_practicals/xschem/7804_AND_IC.sch
.subckt 7804_AND_IC A B Y VCC GND
*.PININFO A:I Y:O B:I VCC:B GND:B
XM2 net1 A VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM3 net1 B VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM5 Y net1 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM1 net1 A net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net2 B GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 Y net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
