** sch_path: /home/iappiah/tt_project2_practicals/xschem/ic_7804_AND.sch
.subckt ic_7804_AND A B Y VCC GND
*.PININFO A:I Y:O B:I VCC:B GND:B
XM2 net1 A VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM3 net1 B VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM5 Y net1 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM1 net1 A net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net2 B GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 Y net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends
.end
