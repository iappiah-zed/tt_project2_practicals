magic
tech sky130A
magscale 1 2
timestamp 1771336497
<< metal1 >>
rect -6124 203 -5924 346
rect -6143 -867 -5900 203
rect -6143 -1110 425 -867
rect 7783 -1110 13707 -867
rect -6143 -13185 -5900 -1110
rect 8862 -2685 9062 -2646
rect -288 -2796 -88 -2748
rect -288 -2905 1075 -2796
rect 7696 -2810 9062 -2685
rect 8862 -2846 9062 -2810
rect 12272 -2689 12472 -2656
rect 12272 -2814 13769 -2689
rect 21382 -2800 21582 -2758
rect 12272 -2856 12472 -2814
rect -288 -2948 -88 -2905
rect 20368 -2909 21582 -2800
rect 21382 -2958 21582 -2909
rect -124 -3810 1126 -3809
rect -288 -4009 1126 -3810
rect 20256 -3814 21378 -3813
rect -288 -4010 -88 -4009
rect 20256 -4013 21574 -3814
rect 21374 -4014 21574 -4013
rect 7855 -5224 13651 -4961
rect 21133 -6917 21396 -4965
rect 21133 -6952 22165 -6917
rect 21133 -7152 22344 -6952
rect 21133 -7180 22165 -7152
rect 7757 -9348 13849 -9085
rect 21133 -9348 21396 -7180
rect -156 -10284 1126 -10282
rect -320 -10482 1126 -10284
rect -320 -10484 -120 -10482
rect 20272 -10496 21584 -10296
rect -324 -11386 -124 -11344
rect -324 -11495 1197 -11386
rect 21384 -11400 21584 -11356
rect 8860 -11481 9060 -11444
rect -324 -11544 -124 -11495
rect 7730 -11606 9060 -11481
rect 8860 -11644 9060 -11606
rect 12270 -11495 12470 -11456
rect 12270 -11620 13669 -11495
rect 20202 -11509 21584 -11400
rect 21384 -11556 21584 -11509
rect 12270 -11656 12470 -11620
rect -6143 -13428 475 -13185
rect 7749 -13442 13609 -13199
use ic_7804_AND  x1
timestamp 1771333935
transform 1 0 599 0 1 -2088
box -587 -3132 7601 1225
use ic_7804_AND  x2
timestamp 1771333935
transform -1 0 20833 0 1 -2092
box -587 -3132 7601 1225
use ic_7804_AND  x3
timestamp 1771333935
transform -1 0 20809 0 -1 -12217
box -587 -3132 7601 1225
use ic_7804_AND  x4
timestamp 1771333935
transform 1 0 577 0 -1 -12203
box -587 -3132 7601 1225
<< labels >>
flabel metal1 -288 -2948 -88 -2748 0 FreeSans 256 0 0 0 1A
port 0 nsew
flabel metal1 -288 -4010 -88 -3810 0 FreeSans 256 0 0 0 1B
port 1 nsew
flabel metal1 8862 -2846 9062 -2646 0 FreeSans 256 0 0 0 1Y
port 2 nsew
flabel metal1 12272 -2856 12472 -2656 0 FreeSans 256 0 0 0 2Y
port 5 nsew
flabel metal1 21382 -2958 21582 -2758 0 FreeSans 256 0 0 0 2A
port 3 nsew
flabel metal1 21374 -4014 21574 -3814 0 FreeSans 256 0 0 0 2B
port 4 nsew
flabel metal1 12270 -11656 12470 -11456 0 FreeSans 256 0 0 0 3Y
port 9 nsew
flabel metal1 21384 -10496 21584 -10296 0 FreeSans 256 0 0 0 3B
port 8 nsew
flabel metal1 21384 -11556 21584 -11356 0 FreeSans 256 0 0 0 3A
port 7 nsew
flabel metal1 8860 -11644 9060 -11444 0 FreeSans 256 0 0 0 4Y
port 12 nsew
flabel metal1 -320 -10484 -120 -10284 0 FreeSans 256 0 0 0 4B
port 11 nsew
flabel metal1 -324 -11544 -124 -11344 0 FreeSans 256 0 0 0 4A
port 10 nsew
flabel metal1 -6124 146 -5924 346 0 FreeSans 256 0 0 0 VCC
port 13 nsew
flabel metal1 22144 -7152 22344 -6952 0 FreeSans 256 0 0 0 GND
port 6 nsew
<< end >>
