** sch_path: /home/iappiah/tt_project2_practicals/xschem/ic_7408_testbench.sch
.subckt ic_7408_testbench 1A GND 1Y 1B 2A 2B 3A 3B 4A 4B 2Y 3Y 4Y VCC
*.PININFO 1A:I GND:B 1Y:O 1B:I 2A:I 2B:I 3A:I 3B:I 4A:I 4B:I 2Y:O 3Y:O 4Y:O VCC:B
V1 VCC GND 1.8
V2 1A GND pulse(0 1.8 1u 1n 1n 2u 4u)
V3 1B GND pulse(0 1.8 1u 1n 1n 2u 4u)
R1 out_1y_before 1Y 1k m=1
C1 1Y GND 10p m=1
x1 1A 1B out_1y_before 2A 2B 2Y GND 3A 3B 3Y 4A 4B 4Y net1 AND_IC_TopLevel
Vmeas VCC net1 0
.save i(vmeas)
R3 out_1y_before1 1Y_out 1k m=1
C3 1Y_out GND 10p m=1
x2 1A 1B out_1y_before1 2A 2B 2Y_out GND 3A 3B 3Y_out 4A 4B 4Y_out net2 AND_IC_TopLevel_parax
Vmeas1 VCC net2 0
.save i(vmeas1)
V4 2A GND 1.8
V5 2B GND 1.8
V6 3A GND 1.8
V7 3B GND 1.8
V8 4A GND 1.8
V9 4B GND 1.8
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/iappiah/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.tran 10n 8u
.save all

.control
run
write 7408IC_final_testbench.raw

.endc



**** end user architecture code
.ends

* expanding   symbol:  AND_IC_TopLevel.sym # of pins=14
** sym_path: /home/iappiah/tt_project2_practicals/xschem/AND_IC_TopLevel.sym
** sch_path: /home/iappiah/tt_project2_practicals/xschem/AND_IC_TopLevel.sch
.subckt AND_IC_TopLevel 1A 1B 1Y 2A 2B 2Y GND 3A 3B 3Y 4A 4B 4Y VCC
*.PININFO 1A:I GND:B 1Y:O 1B:I 2A:I 2B:I 3A:I 3B:I 4A:I 4B:I 2Y:O 3Y:O 4Y:O VCC:B
x1 1A 1B 1Y VCC GND ic_7804_AND
x2 2A 2B 2Y VCC GND ic_7804_AND
x3 3A 3B 3Y VCC GND ic_7804_AND
x4 4A 4B 4Y VCC GND ic_7804_AND
.ends


* expanding   symbol:  AND_IC_TopLevel_parax.sym # of pins=14
** sym_path: /home/iappiah/tt_project2_practicals/xschem/AND_IC_TopLevel.sym
.include /home/iappiah/tt_project2_practicals/mag/AND_IC_TopLevel.sim.spice

* expanding   symbol:  ic_7804_AND.sym # of pins=5
** sym_path: /home/iappiah/tt_project2_practicals/xschem/ic_7804_AND.sym
** sch_path: /home/iappiah/tt_project2_practicals/xschem/ic_7804_AND.sch
.subckt ic_7804_AND A B Y VCC GND
*.PININFO A:I Y:O B:I VCC:B GND:B
XM2 net1 A VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM3 net1 B VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM5 Y net1 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM1 net1 A net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net2 B GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 Y net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.GLOBAL GND
.end
