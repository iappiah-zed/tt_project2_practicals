magic
tech sky130A
magscale 1 2
timestamp 1771524365
<< metal1 >>
rect 1437 33750 1637 33756
rect 1437 33126 1637 33550
rect 6612 31248 6618 31308
rect 6678 31248 6684 31308
rect 7344 31262 7350 31322
rect 7410 31262 7416 31322
rect 6618 29128 6678 31248
rect 7350 30140 7410 31262
rect 16494 31158 16500 31218
rect 16560 31158 16566 31218
rect 16500 30214 16560 31158
rect 19890 31092 19896 31152
rect 19956 31092 19962 31152
rect 19896 30222 19956 31092
rect 28376 30904 28382 30964
rect 28442 30904 28448 30964
rect 28382 30138 28442 30904
rect 28872 29510 28878 29570
rect 28938 29510 28944 29570
rect 6618 29068 7390 29128
rect 28878 29038 28938 29510
rect 29705 25860 30342 26060
rect 28472 23228 28532 23234
rect 28532 23168 29076 23228
rect 28472 23162 28532 23168
rect 6216 22660 6276 22666
rect 6276 22600 7366 22660
rect 6216 22594 6276 22600
rect 29016 22588 29076 23168
rect 16484 22094 16490 22154
rect 16550 22094 16556 22154
rect 19890 22124 19896 22184
rect 19956 22124 19962 22184
rect 6206 21546 6212 21606
rect 6272 21546 7408 21606
rect 16490 21444 16550 22094
rect 19896 21476 19956 22124
rect 29612 21908 29672 21914
rect 29612 21590 29672 21848
rect 29028 21530 29672 21590
rect 30142 21292 30342 25860
rect 30142 21086 30342 21092
<< via1 >>
rect 1437 33550 1637 33750
rect 6618 31248 6678 31308
rect 7350 31262 7410 31322
rect 16500 31158 16560 31218
rect 19896 31092 19956 31152
rect 28382 30904 28442 30964
rect 28878 29510 28938 29570
rect 28472 23168 28532 23228
rect 6216 22600 6276 22660
rect 16490 22094 16550 22154
rect 19896 22124 19956 22184
rect 6212 21546 6272 21606
rect 29612 21848 29672 21908
rect 30142 21092 30342 21292
<< metal2 >>
rect 5644 34210 5704 34212
rect 1437 34164 1637 34173
rect 5637 34154 5646 34210
rect 5702 34154 5711 34210
rect 6618 34206 6678 34208
rect 1437 33750 1637 33964
rect 1431 33550 1437 33750
rect 1637 33550 1643 33750
rect 5644 22660 5704 34154
rect 6611 34150 6620 34206
rect 6676 34150 6685 34206
rect 7352 34204 7408 34211
rect 7350 34202 7410 34204
rect 6618 31308 6678 34150
rect 7350 34146 7352 34202
rect 7408 34146 7410 34202
rect 7350 31322 7410 34146
rect 16500 31362 16560 31364
rect 16493 31306 16502 31362
rect 16558 31306 16567 31362
rect 19896 31334 19956 31336
rect 7350 31256 7410 31262
rect 6618 31242 6678 31248
rect 16500 31218 16560 31306
rect 19889 31278 19898 31334
rect 19954 31278 19963 31334
rect 16500 31152 16560 31158
rect 19896 31152 19956 31278
rect 28382 31254 28442 31256
rect 28375 31198 28384 31254
rect 28440 31198 28449 31254
rect 19896 31086 19956 31092
rect 28382 30964 28442 31198
rect 28382 30898 28442 30904
rect 28878 29706 28938 29708
rect 28871 29650 28880 29706
rect 28936 29650 28945 29706
rect 28878 29570 28938 29650
rect 28878 29504 28938 29510
rect 28050 23228 28106 23235
rect 28048 23226 28472 23228
rect 28048 23170 28050 23226
rect 28106 23170 28472 23226
rect 28048 23168 28472 23170
rect 28532 23168 28538 23228
rect 28050 23161 28106 23168
rect 5644 22600 6216 22660
rect 6276 22600 6282 22660
rect 16490 22490 16550 22492
rect 16483 22434 16492 22490
rect 16548 22434 16557 22490
rect 19896 22470 19956 22472
rect 16490 22154 16550 22434
rect 19889 22414 19898 22470
rect 19954 22414 19963 22470
rect 19896 22184 19956 22414
rect 29612 22166 29672 22168
rect 19896 22118 19956 22124
rect 29605 22110 29614 22166
rect 29670 22110 29679 22166
rect 16490 22088 16550 22094
rect 29612 21908 29672 22110
rect 29606 21848 29612 21908
rect 29672 21848 29678 21908
rect 4568 21606 4624 21613
rect 6212 21606 6272 21612
rect 4566 21604 6212 21606
rect 4566 21548 4568 21604
rect 4624 21548 6212 21604
rect 4566 21546 6212 21548
rect 4568 21539 4624 21546
rect 6212 21540 6272 21546
rect 30136 21092 30142 21292
rect 30342 21092 30348 21292
rect 30142 20230 30342 21092
rect 30142 20021 30342 20030
<< via2 >>
rect 1437 33964 1637 34164
rect 5646 34154 5702 34210
rect 6620 34150 6676 34206
rect 7352 34146 7408 34202
rect 16502 31306 16558 31362
rect 19898 31278 19954 31334
rect 28384 31198 28440 31254
rect 28880 29650 28936 29706
rect 28050 23170 28106 23226
rect 16492 22434 16548 22490
rect 19898 22414 19954 22470
rect 29614 22110 29670 22166
rect 4568 21548 4624 21604
rect 30142 20030 30342 20230
<< metal3 >>
rect 18270 44086 18276 44150
rect 18340 44148 18346 44150
rect 19888 44148 19894 44150
rect 18340 44088 19894 44148
rect 18340 44086 18346 44088
rect 19888 44086 19894 44088
rect 19958 44086 19964 44150
rect 23788 43256 23794 43320
rect 23858 43256 23864 43320
rect 20672 42724 20736 42730
rect 15156 42660 15162 42724
rect 15226 42722 15232 42724
rect 15226 42662 20672 42722
rect 15226 42660 15232 42662
rect 20672 42654 20736 42660
rect 20682 41876 20746 41882
rect 23796 41876 23856 43256
rect 14482 41812 14488 41876
rect 14552 41874 14558 41876
rect 14552 41814 20682 41874
rect 14552 41812 14558 41814
rect 23788 41812 23794 41876
rect 23858 41812 23864 41876
rect 20682 41806 20746 41812
rect 17166 40148 17172 40212
rect 17236 40148 17242 40212
rect 18204 40176 18268 40182
rect 17174 38458 17234 40148
rect 18204 40106 18268 40112
rect 18206 38462 18266 40106
rect 17166 38394 17172 38458
rect 17236 38394 17242 38458
rect 18204 38456 18268 38462
rect 18204 38386 18268 38392
rect 6612 37672 6618 37674
rect 5644 37612 6618 37672
rect 5644 35860 5704 37612
rect 6612 37610 6618 37612
rect 6682 37610 6688 37674
rect 5636 35796 5642 35860
rect 5706 35796 5712 35860
rect 15372 35854 15436 35860
rect 20628 35854 20692 35860
rect 15366 35790 15372 35854
rect 15436 35852 15442 35854
rect 15436 35792 20628 35852
rect 15436 35790 15442 35792
rect 15372 35784 15436 35790
rect 20628 35784 20692 35790
rect 24196 35854 24260 35860
rect 27102 35852 27108 35854
rect 24260 35792 27108 35852
rect 27102 35790 27108 35792
rect 27172 35790 27178 35854
rect 24196 35784 24260 35790
rect 15374 35124 15438 35130
rect 20640 35124 20704 35130
rect 15438 35062 20640 35122
rect 15374 35054 15438 35060
rect 20640 35054 20704 35060
rect 24164 35124 24228 35130
rect 27660 35124 27724 35130
rect 24228 35062 27660 35122
rect 24164 35054 24228 35060
rect 27660 35054 27724 35060
rect 5642 34738 5706 34744
rect 244 34536 250 34736
rect 450 34536 1637 34736
rect 5642 34668 5706 34674
rect 6610 34670 6616 34734
rect 6680 34670 6686 34734
rect 1437 34169 1637 34536
rect 5644 34215 5704 34668
rect 5641 34210 5707 34215
rect 6618 34211 6678 34670
rect 7342 34636 7348 34700
rect 7412 34636 7418 34700
rect 1432 34164 1642 34169
rect 1432 33964 1437 34164
rect 1637 33964 1642 34164
rect 5641 34154 5646 34210
rect 5702 34154 5707 34210
rect 5641 34149 5707 34154
rect 6615 34206 6681 34211
rect 7350 34207 7410 34636
rect 25996 34316 26060 34322
rect 28870 34314 28876 34316
rect 26060 34254 28876 34314
rect 28870 34252 28876 34254
rect 28940 34252 28946 34316
rect 25996 34246 26060 34252
rect 6615 34150 6620 34206
rect 6676 34150 6681 34206
rect 6615 34145 6681 34150
rect 7347 34202 7413 34207
rect 7347 34146 7352 34202
rect 7408 34146 7413 34202
rect 7347 34141 7413 34146
rect 1432 33959 1642 33964
rect 16492 31446 16498 31510
rect 16562 31446 16568 31510
rect 19888 31450 19894 31514
rect 19958 31450 19964 31514
rect 28374 31492 28380 31556
rect 28444 31492 28450 31556
rect 16500 31367 16560 31446
rect 16497 31362 16563 31367
rect 16497 31306 16502 31362
rect 16558 31306 16563 31362
rect 19896 31339 19956 31450
rect 16497 31301 16563 31306
rect 19893 31334 19959 31339
rect 19893 31278 19898 31334
rect 19954 31278 19959 31334
rect 19893 31273 19959 31278
rect 28382 31259 28442 31492
rect 28379 31254 28445 31259
rect 28379 31198 28384 31254
rect 28440 31198 28445 31254
rect 28379 31193 28445 31198
rect 28870 29786 28876 29850
rect 28940 29786 28946 29850
rect 28878 29711 28938 29786
rect 28875 29706 28941 29711
rect 28875 29650 28880 29706
rect 28936 29650 28941 29706
rect 28875 29645 28941 29650
rect 27696 23230 27760 23236
rect 28045 23228 28111 23231
rect 27760 23226 28111 23228
rect 27760 23170 28050 23226
rect 28106 23170 28111 23226
rect 27760 23168 28111 23170
rect 27696 23160 27760 23166
rect 28045 23165 28111 23168
rect 16482 22702 16488 22766
rect 16552 22702 16558 22766
rect 4564 22546 4628 22552
rect 16490 22495 16550 22702
rect 19888 22696 19894 22760
rect 19958 22696 19964 22760
rect 4564 22476 4628 22482
rect 16487 22490 16553 22495
rect 4566 21609 4626 22476
rect 16487 22434 16492 22490
rect 16548 22434 16553 22490
rect 19896 22475 19956 22696
rect 16487 22429 16553 22434
rect 19893 22470 19959 22475
rect 19893 22414 19898 22470
rect 19954 22414 19959 22470
rect 19893 22409 19959 22414
rect 29604 22346 29610 22410
rect 29674 22346 29680 22410
rect 29612 22171 29672 22346
rect 29609 22166 29675 22171
rect 29609 22110 29614 22166
rect 29670 22110 29675 22166
rect 29609 22105 29675 22110
rect 4563 21604 4629 21609
rect 4563 21548 4568 21604
rect 4624 21548 4629 21604
rect 4563 21543 4629 21548
rect 30137 20230 30347 20235
rect 30137 20030 30142 20230
rect 30342 20030 30347 20230
rect 30137 20025 30347 20030
rect 30142 17936 30342 20025
rect 30142 17730 30342 17736
<< via3 >>
rect 18276 44086 18340 44150
rect 19894 44086 19958 44150
rect 23794 43256 23858 43320
rect 15162 42660 15226 42724
rect 20672 42660 20736 42724
rect 14488 41812 14552 41876
rect 20682 41812 20746 41876
rect 23794 41812 23858 41876
rect 17172 40148 17236 40212
rect 18204 40112 18268 40176
rect 17172 38394 17236 38458
rect 18204 38392 18268 38456
rect 6618 37610 6682 37674
rect 5642 35796 5706 35860
rect 15372 35790 15436 35854
rect 20628 35790 20692 35854
rect 24196 35790 24260 35854
rect 27108 35790 27172 35854
rect 15374 35060 15438 35124
rect 20640 35060 20704 35124
rect 24164 35060 24228 35124
rect 27660 35060 27724 35124
rect 250 34536 450 34736
rect 5642 34674 5706 34738
rect 6616 34670 6680 34734
rect 7348 34636 7412 34700
rect 25996 34252 26060 34316
rect 28876 34252 28940 34316
rect 16498 31446 16562 31510
rect 19894 31450 19958 31514
rect 28380 31492 28444 31556
rect 28876 29786 28940 29850
rect 27696 23166 27760 23230
rect 16488 22702 16552 22766
rect 4564 22482 4628 22546
rect 19894 22696 19958 22760
rect 29610 22346 29674 22410
rect 30142 17736 30342 17936
<< metal4 >>
rect 6134 44754 6194 45152
rect 6686 44754 6746 45152
rect 7238 44754 7298 45152
rect 7790 44754 7850 45152
rect 8342 44754 8402 45152
rect 8894 44754 8954 45152
rect 9446 44754 9506 45152
rect 9998 44754 10058 45152
rect 10550 44754 10610 45152
rect 11102 44754 11162 45152
rect 11654 44754 11714 45152
rect 12206 44754 12266 45152
rect 12758 44754 12818 45152
rect 13310 44754 13370 45152
rect 13862 44754 13922 45152
rect 14414 44754 14474 45152
rect 14966 44754 15026 45152
rect 15518 44754 15578 45152
rect 16070 44754 16130 45152
rect 16622 44754 16682 45152
rect 6118 44674 16682 44754
rect 6118 44672 16673 44674
rect 200 34736 600 44152
rect 200 34536 250 34736
rect 450 34536 600 34736
rect 200 1000 600 34536
rect 800 43971 1200 44152
rect 6118 43971 6200 44672
rect 8894 44670 8954 44672
rect 14414 44670 14474 44672
rect 800 43889 6200 43971
rect 800 18026 1200 43889
rect 15161 42724 15227 42725
rect 15161 42660 15162 42724
rect 15226 42660 15227 42724
rect 15161 42659 15227 42660
rect 14487 41876 14553 41877
rect 14487 41812 14488 41876
rect 14552 41812 14553 41876
rect 14487 41811 14553 41812
rect 6617 37674 6683 37675
rect 6617 37610 6618 37674
rect 6682 37672 6683 37674
rect 14490 37672 14550 41811
rect 6682 37612 14550 37672
rect 6682 37610 6683 37612
rect 6617 37609 6683 37610
rect 15164 36756 15224 42659
rect 17174 40213 17234 45152
rect 17726 41092 17786 45152
rect 18278 44151 18338 45152
rect 18275 44150 18341 44151
rect 18275 44086 18276 44150
rect 18340 44086 18341 44150
rect 18275 44085 18341 44086
rect 17726 41032 18266 41092
rect 17171 40212 17237 40213
rect 17171 40148 17172 40212
rect 17236 40148 17237 40212
rect 18206 40177 18266 41032
rect 17171 40147 17237 40148
rect 18203 40176 18269 40177
rect 18203 40112 18204 40176
rect 18268 40112 18269 40176
rect 18203 40111 18269 40112
rect 18830 39256 18890 45152
rect 19382 44950 19442 45152
rect 19934 44950 19994 45152
rect 20486 44950 20546 45152
rect 21038 44950 21098 45152
rect 21590 44950 21650 45152
rect 22142 44950 22202 45152
rect 22694 44950 22754 45152
rect 23246 44950 23306 45152
rect 23798 44582 23858 45152
rect 23796 44454 23858 44582
rect 19893 44150 19959 44151
rect 19893 44086 19894 44150
rect 19958 44086 19959 44150
rect 19893 44085 19959 44086
rect 4566 36696 15224 36756
rect 16500 39196 18890 39256
rect 4566 22547 4626 36696
rect 5641 35860 5707 35861
rect 5641 35796 5642 35860
rect 5706 35796 5707 35860
rect 15371 35854 15437 35855
rect 15371 35852 15372 35854
rect 5641 35795 5707 35796
rect 5644 34739 5704 35795
rect 6618 35792 15372 35852
rect 5641 34738 5707 34739
rect 5641 34674 5642 34738
rect 5706 34674 5707 34738
rect 6618 34735 6678 35792
rect 15371 35790 15372 35792
rect 15436 35790 15437 35854
rect 15371 35789 15437 35790
rect 15373 35124 15439 35125
rect 15373 35122 15374 35124
rect 7350 35062 15374 35122
rect 5641 34673 5707 34674
rect 6615 34734 6681 34735
rect 6615 34670 6616 34734
rect 6680 34670 6681 34734
rect 7350 34701 7410 35062
rect 15373 35060 15374 35062
rect 15438 35060 15439 35124
rect 15373 35059 15439 35060
rect 6615 34669 6681 34670
rect 7347 34700 7413 34701
rect 7347 34636 7348 34700
rect 7412 34636 7413 34700
rect 7347 34635 7413 34636
rect 16500 31511 16560 39196
rect 17171 38458 17237 38459
rect 17171 38394 17172 38458
rect 17236 38394 17237 38458
rect 17171 38393 17237 38394
rect 18203 38456 18269 38457
rect 16497 31510 16563 31511
rect 16497 31446 16498 31510
rect 16562 31446 16563 31510
rect 16497 31445 16563 31446
rect 17174 23064 17234 38393
rect 18203 38392 18204 38456
rect 18268 38454 18269 38456
rect 18268 38394 18886 38454
rect 18268 38392 18269 38394
rect 18203 38391 18269 38392
rect 16490 23004 17234 23064
rect 18826 23064 18886 38394
rect 19896 31515 19956 44085
rect 23796 43321 23856 44454
rect 24350 44364 24410 45152
rect 24348 44222 24410 44364
rect 23793 43320 23859 43321
rect 23793 43256 23794 43320
rect 23858 43256 23859 43320
rect 23793 43255 23859 43256
rect 20671 42724 20737 42725
rect 20671 42660 20672 42724
rect 20736 42722 20737 42724
rect 24348 42722 24408 44222
rect 20736 42662 24408 42722
rect 20736 42660 20737 42662
rect 20671 42659 20737 42660
rect 20681 41876 20747 41877
rect 20681 41812 20682 41876
rect 20746 41874 20747 41876
rect 23793 41876 23859 41877
rect 23793 41874 23794 41876
rect 20746 41814 23794 41874
rect 20746 41812 20747 41814
rect 20681 41811 20747 41812
rect 23793 41812 23794 41814
rect 23858 41812 23859 41876
rect 23793 41811 23859 41812
rect 20627 35854 20693 35855
rect 20627 35790 20628 35854
rect 20692 35852 20693 35854
rect 24195 35854 24261 35855
rect 24195 35852 24196 35854
rect 20692 35792 24196 35852
rect 20692 35790 20693 35792
rect 20627 35789 20693 35790
rect 24195 35790 24196 35792
rect 24260 35790 24261 35854
rect 24195 35789 24261 35790
rect 20639 35124 20705 35125
rect 20639 35060 20640 35124
rect 20704 35122 20705 35124
rect 24163 35124 24229 35125
rect 24163 35122 24164 35124
rect 20704 35062 24164 35122
rect 20704 35060 20705 35062
rect 20639 35059 20705 35060
rect 24163 35060 24164 35062
rect 24228 35060 24229 35124
rect 24163 35059 24229 35060
rect 24902 33534 24962 45152
rect 20974 33474 24962 33534
rect 19893 31514 19959 31515
rect 19893 31450 19894 31514
rect 19958 31450 19959 31514
rect 19893 31449 19959 31450
rect 20974 26336 21034 33474
rect 25454 32914 25514 45152
rect 26006 44463 26066 45152
rect 25985 41003 26071 44463
rect 25998 34317 26058 41003
rect 25995 34316 26061 34317
rect 25995 34252 25996 34316
rect 26060 34252 26061 34316
rect 25995 34251 26061 34252
rect 23994 32854 25514 32914
rect 26558 32894 26618 45152
rect 27110 35855 27170 45152
rect 27107 35854 27173 35855
rect 27107 35790 27108 35854
rect 27172 35790 27173 35854
rect 27107 35789 27173 35790
rect 27662 35125 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27659 35124 27725 35125
rect 27659 35060 27660 35124
rect 27724 35060 27725 35124
rect 27659 35059 27725 35060
rect 28875 34316 28941 34317
rect 28875 34252 28876 34316
rect 28940 34252 28941 34316
rect 28875 34251 28941 34252
rect 23994 26902 24054 32854
rect 26558 32834 28442 32894
rect 28382 31557 28442 32834
rect 28379 31556 28445 31557
rect 28379 31492 28380 31556
rect 28444 31492 28445 31556
rect 28379 31491 28445 31492
rect 28878 29851 28938 34251
rect 28875 29850 28941 29851
rect 28875 29786 28876 29850
rect 28940 29786 28941 29850
rect 28875 29785 28941 29786
rect 23994 26842 28054 26902
rect 20974 26276 27398 26336
rect 27338 23228 27398 26276
rect 27994 25234 28054 26842
rect 27994 25174 29672 25234
rect 27695 23230 27761 23231
rect 27695 23228 27696 23230
rect 27338 23168 27696 23228
rect 27695 23166 27696 23168
rect 27760 23166 27761 23230
rect 27695 23165 27761 23166
rect 18826 23004 19956 23064
rect 16490 22767 16550 23004
rect 16487 22766 16553 22767
rect 16487 22702 16488 22766
rect 16552 22702 16553 22766
rect 19896 22761 19956 23004
rect 16487 22701 16553 22702
rect 19893 22760 19959 22761
rect 19893 22696 19894 22760
rect 19958 22696 19959 22760
rect 19893 22695 19959 22696
rect 4563 22546 4629 22547
rect 4563 22482 4564 22546
rect 4628 22482 4629 22546
rect 4563 22481 4629 22482
rect 29612 22411 29672 25174
rect 29609 22410 29675 22411
rect 29609 22346 29610 22410
rect 29674 22346 29675 22410
rect 29609 22345 29675 22346
rect 800 17936 29072 18026
rect 30141 17936 30343 17937
rect 800 17736 30142 17936
rect 30342 17736 30343 17936
rect 800 17626 29072 17736
rect 30141 17735 30343 17736
rect 800 1000 1200 17626
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use AND_IC_TopLevel  AND_IC_TopLevel_0
timestamp 1771336497
transform 1 0 7561 0 1 33012
box -6143 -13442 22344 346
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
