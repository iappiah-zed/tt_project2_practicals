magic
tech sky130A
magscale 1 2
timestamp 1771244448
<< viali >>
rect 5056 14522 5134 14576
rect 12395 14539 12471 14587
rect 31368 14586 31436 14636
rect 24084 14518 24162 14566
rect 5052 13982 5138 14028
rect 12396 14006 12466 14054
rect 31366 14046 31438 14094
rect 24080 13984 24158 14030
rect 5086 12066 5156 12112
rect 31386 12044 31456 12094
rect 5080 11482 5154 11528
rect 31376 11486 31464 11532
rect 1546 10632 1618 10678
rect 31256 1584 31304 1660
rect 5122 1496 5170 1570
rect 31376 1090 31446 1142
rect 4978 900 5048 948
rect 4978 -582 5054 -534
rect 13212 -544 13286 -498
rect 24090 -552 24160 -504
rect 31262 -802 31308 -732
rect 4986 -1206 5056 -1156
rect 13212 -1174 13282 -1124
rect 24090 -1172 24162 -1120
rect 31384 -1288 31454 -1236
<< metal1 >>
rect 2335 15350 5268 15357
rect 546 15114 5268 15350
rect 546 15106 2910 15114
rect 546 10826 790 15106
rect 3861 14939 3951 15114
rect 3855 14849 3861 14939
rect 3951 14849 3957 14939
rect 5056 14642 5138 15114
rect 12388 14646 12478 15221
rect 12551 15144 23959 15387
rect 12623 15114 12872 15144
rect 24068 14622 24174 15212
rect 5046 14576 5150 14596
rect 5046 14522 5056 14576
rect 5134 14522 5150 14576
rect 5046 14449 5150 14522
rect 12379 14587 12485 14595
rect 12379 14539 12395 14587
rect 12471 14539 12485 14587
rect 12379 14466 12485 14539
rect 4646 14345 5150 14449
rect 3861 14335 3951 14341
rect 1852 13407 2052 13452
rect 3194 13407 3303 13413
rect 1852 13298 3194 13407
rect 1852 13252 2052 13298
rect 3194 13292 3303 13298
rect 1846 12720 2046 12744
rect 1846 12592 3214 12720
rect 3342 12592 3348 12720
rect 1846 12544 2046 12592
rect 3861 12266 3951 14245
rect 4646 13407 4750 14345
rect 5046 14089 5150 14345
rect 12018 14360 12485 14466
rect 5038 14028 5152 14042
rect 5038 13982 5052 14028
rect 5138 13982 5152 14028
rect 5038 13675 5152 13982
rect 5038 13555 5152 13561
rect 6558 13469 6602 13539
rect 5542 13422 6602 13469
rect 12018 13424 12124 14360
rect 12379 14097 12485 14360
rect 24064 14566 24176 14574
rect 24064 14518 24084 14566
rect 24162 14518 24176 14566
rect 24064 14458 24176 14518
rect 24064 14346 24512 14458
rect 24064 14092 24176 14346
rect 12376 14054 12486 14062
rect 12376 14006 12396 14054
rect 12466 14006 12486 14054
rect 12376 13926 12486 14006
rect 24060 14030 24182 14042
rect 24060 13984 24080 14030
rect 24158 13984 24182 14030
rect 24060 13952 24182 13984
rect 12376 13810 12486 13816
rect 24062 13863 24180 13952
rect 24062 13739 24180 13745
rect 5464 13414 6602 13422
rect 5464 13407 6566 13414
rect 4170 13298 4176 13407
rect 4285 13298 6566 13407
rect 12762 13374 13972 13574
rect 22682 13565 22882 13602
rect 22682 13440 24082 13565
rect 24400 13468 24512 14346
rect 29614 14102 29678 15188
rect 31348 14690 31458 15192
rect 31346 14636 31460 14644
rect 31346 14586 31368 14636
rect 31436 14586 31460 14636
rect 31346 14517 31460 14586
rect 31346 14403 31857 14517
rect 31346 14154 31460 14403
rect 29608 14038 29614 14102
rect 29678 14038 29684 14102
rect 31344 14094 31460 14100
rect 31344 14046 31366 14094
rect 31438 14046 31460 14094
rect 31344 13966 31458 14046
rect 30992 13636 30998 13688
rect 31050 13683 31056 13688
rect 31383 13683 31425 13966
rect 31050 13641 31425 13683
rect 31050 13636 31056 13641
rect 31743 13454 31857 14403
rect 32436 13454 32636 13496
rect 22682 13402 22882 13440
rect 30719 13345 32636 13454
rect 5542 13274 6566 13298
rect 5464 13269 6566 13274
rect 24056 13201 24062 13319
rect 24180 13201 24186 13319
rect 32436 13296 32636 13345
rect 12370 12953 12376 13063
rect 12486 12953 12492 13063
rect 4214 12592 4220 12720
rect 4348 12592 5601 12720
rect 3861 12176 5168 12266
rect 5473 12255 5601 12592
rect 5066 12112 5170 12124
rect 5066 12066 5086 12112
rect 5156 12066 5170 12112
rect 4417 11997 4531 12003
rect 4417 11263 4531 11883
rect 5066 11980 5170 12066
rect 5480 11980 5584 12255
rect 5066 11876 5584 11980
rect 5066 11584 5170 11876
rect 5058 11528 5176 11537
rect 5058 11482 5080 11528
rect 5154 11482 5176 11528
rect 5058 11263 5176 11482
rect 12376 11263 12486 12953
rect 17700 11263 18084 11266
rect 2335 11000 5220 11263
rect 12376 11067 23919 11263
rect 24062 11101 24180 13201
rect 30400 13134 30464 13140
rect 30400 13022 30464 13070
rect 30400 12958 31468 13022
rect 31374 12893 31468 12958
rect 31368 12799 31374 12893
rect 31468 12799 31474 12893
rect 30049 12763 30127 12769
rect 32434 12734 32634 12762
rect 12454 11000 23919 11067
rect 30049 11053 30127 12685
rect 30905 12606 32634 12734
rect 30905 12314 31036 12606
rect 31374 12475 31468 12481
rect 30905 12277 30917 12314
rect 31027 12277 31033 12314
rect 31374 12152 31468 12381
rect 31366 12094 31476 12100
rect 31366 12044 31386 12094
rect 31456 12044 31476 12094
rect 31366 11979 31476 12044
rect 31741 11979 31851 12606
rect 32434 12562 32634 12606
rect 31366 11869 31851 11979
rect 31366 11594 31476 11869
rect 31364 11532 31478 11540
rect 31364 11486 31376 11532
rect 31464 11486 31478 11532
rect 31364 11163 31478 11486
rect 546 10738 1628 10826
rect 546 -1807 790 10738
rect 1526 10678 1638 10694
rect 1526 10632 1546 10678
rect 1618 10632 1638 10678
rect 1526 2228 1638 10632
rect 17700 2307 18084 11000
rect 2973 2231 5486 2307
rect 2973 2228 5583 2231
rect 1526 2116 5583 2228
rect 2973 2044 5583 2116
rect 5477 1586 5583 2044
rect 4955 1256 5073 1575
rect 5114 1570 5583 1586
rect 5114 1496 5122 1570
rect 5170 1496 5583 1570
rect 5114 1480 5583 1496
rect 4955 1138 5624 1256
rect 4955 948 5073 1138
rect 4955 900 4978 948
rect 5048 900 5073 948
rect 4955 891 5073 900
rect 5506 844 5624 1138
rect 3795 838 3881 844
rect 3881 752 5062 838
rect 3795 746 3881 752
rect 1852 528 2052 570
rect 5506 528 5623 844
rect 6433 661 6539 2183
rect 6433 549 6539 555
rect 1852 411 5623 528
rect 12152 426 12268 2222
rect 12502 2202 24095 2307
rect 12502 2044 24178 2202
rect 17700 2030 18084 2044
rect 24074 1716 24178 2044
rect 24068 1612 24074 1716
rect 24178 1612 24184 1716
rect 30020 630 30085 2206
rect 30916 1674 31024 2204
rect 30916 1660 31314 1674
rect 30916 1584 31256 1660
rect 31304 1584 31314 1660
rect 30916 1566 31314 1584
rect 31352 1365 31466 1668
rect 31352 1251 31923 1365
rect 31352 1142 31466 1251
rect 31352 1090 31376 1142
rect 31446 1090 31466 1142
rect 31352 1074 31466 1090
rect 30020 559 30085 565
rect 30872 586 31004 1066
rect 31356 748 31464 1026
rect 31356 746 31374 748
rect 31446 746 31464 748
rect 31374 670 31446 676
rect 31809 586 31923 1251
rect 32428 586 32628 618
rect 30872 454 32628 586
rect 1852 370 2052 411
rect 12152 310 13308 426
rect 32428 418 32628 454
rect 1850 -6 2050 32
rect 1850 -115 5655 -6
rect 1850 -126 4674 -115
rect 1850 -168 2050 -126
rect 3795 -419 3881 -413
rect 3795 -1807 3881 -505
rect 4554 -934 4674 -126
rect 12590 -228 12973 -103
rect 13098 -228 13104 -103
rect 5857 -323 5963 -317
rect 4964 -429 5857 -323
rect 4964 -534 5070 -429
rect 5857 -435 5963 -429
rect 4964 -582 4978 -534
rect 5054 -582 5070 -534
rect 4964 -594 5070 -582
rect 4956 -934 5076 -648
rect 4554 -1054 5076 -934
rect 12800 -896 12924 -228
rect 13192 -498 13308 310
rect 30798 288 30870 294
rect 29650 216 29656 288
rect 29728 216 30798 288
rect 30798 210 30870 216
rect 32430 -4 32630 38
rect 13405 -103 13530 -97
rect 13738 -103 13938 -66
rect 13530 -228 13938 -103
rect 13405 -234 13530 -228
rect 13738 -266 13938 -228
rect 22702 -99 22902 -60
rect 22702 -224 23931 -99
rect 30699 -113 32630 -4
rect 22702 -260 22902 -224
rect 13192 -544 13212 -498
rect 13286 -544 13308 -498
rect 13192 -546 13308 -544
rect 13194 -556 13308 -546
rect 24074 -358 24178 -352
rect 24074 -504 24178 -462
rect 24074 -552 24090 -504
rect 24160 -552 24178 -504
rect 24074 -564 24178 -552
rect 13186 -896 13310 -612
rect 12800 -1020 13310 -896
rect 4956 -1156 5076 -1054
rect 4956 -1206 4986 -1156
rect 5056 -1206 5076 -1156
rect 13186 -1124 13310 -1020
rect 13186 -1174 13212 -1124
rect 13282 -1174 13310 -1124
rect 13186 -1188 13310 -1174
rect 24068 -907 24182 -618
rect 24375 -907 24489 -121
rect 30558 -330 30623 -324
rect 30623 -395 31047 -330
rect 30558 -401 30623 -395
rect 24068 -1021 24489 -907
rect 29656 -616 29728 -610
rect 24068 -1120 24182 -1021
rect 24068 -1172 24090 -1120
rect 24162 -1172 24182 -1120
rect 24068 -1188 24182 -1172
rect 4956 -1226 5076 -1206
rect 4976 -1354 5497 -1268
rect 546 -2050 5395 -1807
rect 5411 -1977 5497 -1354
rect 12228 -1320 13292 -1240
rect 12228 -1994 12308 -1320
rect 12415 -2046 24049 -1803
rect 24076 -1984 24176 -1238
rect 29656 -2026 29728 -688
rect 30982 -735 31047 -395
rect 31264 -714 31314 -712
rect 31162 -732 31320 -714
rect 31162 -735 31262 -732
rect 30982 -800 31262 -735
rect 31162 -802 31262 -800
rect 31308 -802 31320 -732
rect 31162 -822 31320 -802
rect 31356 -1022 31474 -726
rect 31804 -1022 31920 -113
rect 32430 -162 32630 -113
rect 31356 -1138 31920 -1022
rect 31356 -1236 31474 -1138
rect 31356 -1288 31384 -1236
rect 31454 -1288 31474 -1236
rect 31356 -1296 31474 -1288
rect 31376 -1969 31458 -1354
rect 546 -2072 790 -2050
<< via1 >>
rect 3861 14849 3951 14939
rect 3861 14245 3951 14335
rect 3194 13298 3303 13407
rect 3214 12592 3342 12720
rect 5038 13561 5152 13675
rect 12376 13816 12486 13926
rect 24062 13745 24180 13863
rect 4176 13298 4285 13407
rect 29614 14038 29678 14102
rect 30998 13636 31050 13688
rect 24062 13201 24180 13319
rect 12376 12953 12486 13063
rect 4220 12592 4348 12720
rect 4417 11883 4531 11997
rect 30400 13070 30464 13134
rect 31374 12799 31468 12893
rect 30049 12685 30127 12763
rect 31374 12381 31468 12475
rect 3795 752 3881 838
rect 6433 555 6539 661
rect 24074 1612 24178 1716
rect 30020 565 30085 630
rect 31374 676 31446 748
rect 3795 -505 3881 -419
rect 12973 -228 13098 -103
rect 5857 -429 5963 -323
rect 29656 216 29728 288
rect 30798 216 30870 288
rect 13405 -228 13530 -103
rect 24074 -462 24178 -358
rect 30558 -395 30623 -330
rect 29656 -688 29728 -616
<< metal2 >>
rect 3861 14939 3951 14945
rect 3861 14335 3951 14849
rect 3855 14245 3861 14335
rect 3951 14245 3957 14335
rect 29614 14102 29678 14108
rect 12370 13816 12376 13926
rect 12486 13816 12492 13926
rect 4417 13561 5038 13675
rect 5152 13561 5158 13675
rect 4176 13407 4285 13413
rect 3188 13298 3194 13407
rect 3303 13298 4176 13407
rect 4176 13292 4285 13298
rect 3214 12720 3342 12726
rect 4220 12720 4348 12726
rect 3342 12592 4220 12720
rect 3214 12586 3342 12592
rect 4220 12586 4348 12592
rect 4417 11997 4531 13561
rect 12376 13063 12486 13816
rect 24056 13745 24062 13863
rect 24180 13745 24186 13863
rect 24062 13319 24180 13745
rect 29614 13658 29678 14038
rect 30998 13688 31050 13694
rect 30677 13683 30755 13684
rect 29614 13594 30464 13658
rect 24062 13195 24180 13201
rect 30400 13134 30464 13594
rect 30677 13641 30998 13683
rect 30394 13070 30400 13134
rect 30464 13070 30470 13134
rect 12376 12947 12486 12953
rect 30677 12901 30755 13641
rect 30998 13630 31050 13636
rect 30049 12823 30755 12901
rect 31374 12893 31468 12899
rect 30049 12763 30127 12823
rect 30043 12685 30049 12763
rect 30127 12685 30133 12763
rect 31374 12475 31468 12799
rect 31368 12381 31374 12475
rect 31468 12381 31474 12475
rect 4411 11883 4417 11997
rect 4531 11883 4537 11997
rect 24074 1716 24178 1722
rect 3789 752 3795 838
rect 3881 752 3887 838
rect 3795 -419 3881 752
rect 6427 555 6433 661
rect 6539 555 6545 661
rect 6433 373 6539 555
rect 5857 267 6539 373
rect 5857 -323 5963 267
rect 12973 -103 13098 -97
rect 13098 -228 13405 -103
rect 13530 -228 13536 -103
rect 12973 -234 13098 -228
rect 3789 -505 3795 -419
rect 3881 -505 3887 -419
rect 5851 -429 5857 -323
rect 5963 -429 5969 -323
rect 24074 -358 24178 1612
rect 31368 676 31374 748
rect 31446 676 31452 748
rect 30014 565 30020 630
rect 30085 565 30623 630
rect 29656 288 29728 294
rect 24068 -462 24074 -358
rect 24178 -462 24184 -358
rect 29656 -616 29728 216
rect 30558 -330 30623 565
rect 31374 288 31446 676
rect 30792 216 30798 288
rect 30870 216 31446 288
rect 30552 -395 30558 -330
rect 30623 -395 30629 -330
rect 29650 -688 29656 -616
rect 29728 -688 29734 -616
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D1
timestamp 1770916899
transform 1 0 5097 0 1 14681
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D2
timestamp 1770916899
transform 1 0 5095 0 1 14135
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D3
timestamp 1770916899
transform 1 0 5121 0 1 12219
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D4
timestamp 1770916899
transform 1 0 5117 0 1 11637
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D5
timestamp 1770916899
transform 1 0 12435 0 1 14693
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D6
timestamp 1770916899
transform 1 0 12431 0 1 14161
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D7
timestamp 1770916899
transform 1 0 24121 0 1 14671
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D8
timestamp 1770916899
transform 1 0 24121 0 1 14137
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D9
timestamp 1770916899
transform 1 0 31421 0 1 12199
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D10
timestamp 1770916899
transform 1 0 31421 0 1 11641
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D11
timestamp 1770916899
transform 1 0 31403 0 1 14741
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D12
timestamp 1770916899
transform 1 0 31403 0 1 14201
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D13
timestamp 1770916899
transform 1 0 5017 0 1 795
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D14
timestamp 1770916899
transform 1 0 5015 0 1 1533
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D15
timestamp 1770916899
transform 1 0 5019 0 1 -1311
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D16
timestamp 1770916899
transform 1 0 5017 0 1 -689
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D17
timestamp 1770916899
transform 1 0 31417 0 1 -1391
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D18
timestamp 1770916899
transform 1 0 31417 0 1 -767
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D19
timestamp 1770916899
transform 1 0 31411 0 1 985
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D20
timestamp 1770916899
transform 1 0 31411 0 1 1621
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D21
timestamp 1770916899
transform 1 0 13247 0 1 -1279
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D22
timestamp 1770916899
transform 1 0 13249 0 1 -651
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D23
timestamp 1770916899
transform 1 0 24125 0 1 -1277
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D24
timestamp 1770916899
transform 1 0 24125 0 1 -657
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D25
timestamp 1770916899
transform 1 0 1583 0 1 10783
box -183 -183 183 183
use 7804_AND_IC  x1
timestamp 1770916899
transform 1 0 5361 0 1 14132
box -587 -3132 7601 1225
use 7804_AND_IC  x2
timestamp 1770916899
transform -1 0 31173 0 1 14162
box -587 -3132 7601 1225
use 7804_AND_IC  x3
timestamp 1770916899
transform -1 0 31149 0 -1 -821
box -587 -3132 7601 1225
use 7804_AND_IC  x4
timestamp 1770916899
transform 1 0 5357 0 -1 -825
box -587 -3132 7601 1225
<< labels >>
flabel metal1 1852 13252 2052 13452 0 FreeSans 256 0 0 0 1A
port 0 nsew
flabel metal1 1846 12544 2046 12744 0 FreeSans 256 0 0 0 1B
port 1 nsew
flabel metal1 32436 13296 32636 13496 0 FreeSans 256 0 0 0 2A
port 3 nsew
flabel metal1 32434 12562 32634 12762 0 FreeSans 256 0 0 0 2B
port 4 nsew
flabel metal1 22682 13402 22882 13602 0 FreeSans 256 0 0 0 2Y
port 5 nsew
flabel metal1 13772 13374 13972 13574 0 FreeSans 256 0 0 0 1Y
port 2 nsew
flabel metal1 32430 -162 32630 38 0 FreeSans 256 0 0 0 3A
port 7 nsew
flabel metal1 32428 418 32628 618 0 FreeSans 256 0 0 0 3B
port 8 nsew
flabel metal1 22702 -260 22902 -60 0 FreeSans 256 0 0 0 3Y
port 9 nsew
flabel metal1 13738 -266 13938 -66 0 FreeSans 256 0 0 0 4Y
port 12 nsew
flabel metal1 1850 -168 2050 32 0 FreeSans 256 0 0 0 4A
port 10 nsew
flabel metal1 1852 370 2052 570 0 FreeSans 256 0 0 0 4B
port 11 nsew
flabel metal1 17800 7120 18000 7320 0 FreeSans 256 0 0 0 GND
port 6 nsew
flabel metal1 570 7456 770 7656 0 FreeSans 256 0 0 0 VCC
port 13 nsew
<< end >>
